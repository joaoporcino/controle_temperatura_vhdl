library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top_level is
    Port (
        clk_50MHz : in  STD_LOGIC;
        rst       : in  STD_LOGIC;
        
        -- Entradas
        temp_int_min : in STD_LOGIC_VECTOR(6 downto 0);
        temp_ext_max : in STD_LOGIC_VECTOR(6 downto 0);

        -- Saídas Visuais (LEDs de Estado)
        led_heat   : out STD_LOGIC;
        led_cool   : out STD_LOGIC;
        led_stable : out STD_LOGIC;
        led_alert  : out STD_LOGIC;
        
        motor_pow_c : out STD_LOGIC; -- Sinal de força para Resfriar
        motor_pow_h : out STD_LOGIC; -- Sinal de força para Aquecer
        
        -- Saída de Dados
        power_out  : out STD_LOGIC_VECTOR(6 downto 0);
        
        -- Displays
        hex0       : out STD_LOGIC_VECTOR(6 downto 0);
        hex1       : out STD_LOGIC_VECTOR(6 downto 0)
    );
end top_level;

architecture Structural of top_level is

    component clock_divider is
        Port ( clk_in : in STD_LOGIC; rst : in STD_LOGIC; clk_out : out STD_LOGIC );
    end component;

    component control_decoder is
        Port ( reset : in STD_LOGIC; not_reset : out STD_LOGIC );
    end component;

    signal clk_sys : STD_LOGIC; 

    -- Fios de Controle
    signal w_enab_max, w_enab_min : STD_LOGIC;
    signal w_enab_ext, w_enab_int : STD_LOGIC;
    signal w_enab_pow, w_enab_flags : STD_LOGIC;
    signal control_sw : STD_LOGIC;

    -- Fios de Flags
    signal w_flag_c, w_flag_h, w_flag_s : STD_LOGIC;

begin

    -- Inversor de Reset para Control
    -- Quando rst = '1' (ativo), control_sw = '0' (sistema parado)
    -- Quando rst = '0' (inativo), control_sw = '1' (sistema rodando)
    U_CONTROL_DEC: control_decoder
        port map ( reset => rst, not_reset => control_sw );

    U_CLK_DIV: clock_divider
        port map ( clk_in => clk_50MHz, rst => rst, clk_out => clk_sys );

    U_CONTROLLER: entity work.controller
        port map (
            clk        => clk_sys,
            rst        => rst,
            control    => control_sw,
            c          => w_flag_c,
            h          => w_flag_h,
            s          => w_flag_s,
            enab_max   => w_enab_max,
            enab_min   => w_enab_min,
            enab_ext   => w_enab_ext,
            enab_int   => w_enab_int,
            enab_pow   => w_enab_pow,
            enab_flags => w_enab_flags, 
            heat_out   => led_heat,
            cool_out   => led_cool,
            stable_out => led_stable
        );

    U_DATAPATH: entity work.datapath
        port map (
            clk          => clk_sys,
            rst          => rst,
            temp_int_min => temp_int_min,
            temp_ext_max => temp_ext_max,
            enab_max     => w_enab_max,
            enab_min     => w_enab_min,
            enab_ext     => w_enab_ext,
            enab_int     => w_enab_int,
            enab_pow     => w_enab_pow,
            enab_flags   => w_enab_flags,
            c            => w_flag_c,
            h            => w_flag_h,
            s            => w_flag_s,

            pow_c        => motor_pow_c, 
            pow_h        => motor_pow_h,
            
            alert        => led_alert,
            power_out    => power_out,
            hex0         => hex0,
            hex1         => hex1
        );

end Structural;